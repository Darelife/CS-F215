module mod10_counter (
    input wire clk,
    input wire rst,
    output reg [3:0] count
);
   
    
endmodule