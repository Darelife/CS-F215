`include "dff.v"

module mod16_counter (
    input wire clk,   
    input wire rst,   
    output wire [3:0] q  
);



endmodule
