module preg (
  input clk,
  input reset,
  input [3:0] I,
  output [3:0] A
);
  
endmodule